`timescale 1ns / 1ps
module BitwiseG(
	input Ai,
	input Bi,
	output Gi
    );

and #0.1 (Gi,Ai,Bi);

endmodule
