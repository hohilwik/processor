`timescale 1ns/ 1ps

module fetch_ins(clk, PC, icode, ifun, rA, rB, valC, valP, instr_validity, imem_error, hlt, proc_mem); //(
	input clk;
	input [63:0] PC;
	output reg [3:0] icode;
	output reg [3:0] ifun;
	output reg [3:0] rA;
	output reg [3:0] rB;
	output reg [63:0] valC;
	output reg [63:0] valP;
	output reg instr_validity;
	output reg imem_error;
	output reg hlt;
	output reg [7:0] proc_mem[0:4095];
	//};
	
	//reg [7:0] proc_mem[0:4095];
	reg [0:79] instr; // max instruction length is 10 bytes
	reg [79:0] instr2;
	
	// placeholder for scanf simplicity
	reg [0:7] buffer[0:4095];
	
	
	integer asm_bin_p; // file pointer for binary file
	integer iterlines=0, iterbits=0;
	integer ii=0;
	integer status;
	reg tempbit;
	
	//integer index;
	//initial $readmemb("prog_binary.out",proc_mem);
	//always @index DATA_REG = memory[index];
	
	initial begin
		//$display("%x", buffer[0]);
	   // read from binary file and load into memory
	   
	   //$readmemb("prog_binary.out", buffer);
	   //while(ii<20)
	   //begin
		//$display("%8b", buffer[ii]);
		//ii = ii+1;
	   //end
	   //while(ii<190)
	   //begin
		//  proc_mem[ii] = buffer[ii];
	   //end
	   
	   //asm_bin_p = $fopen("prog_binary.out", "r");
	   //while( !$feof(asm_bin_p) ) 
	   //begin
			
			//status = $fscanf(asm_bin_p, "%b", buffer[0]);
			//$display("%b", buffer[0]);
			//proc_mem[ii] = buffer[0];
			//ii = ii+1;
			//proc_mem[ii] = buffer[ii];
			//ii = ii+1;
			//$fscanf(asm_bin_p, "%b", tempbit);
			//buffer[iterlines][iterbits] = tempbit;
			//iterbits=iterbits+1;
			//if(iterbits>=8) 
			//begin
			//	iterlines=iterlines+1;
			//	iterbits=0;
			//end
				
		//end
		//while(ii<=2000)
		//begin
		//	proc_mem[ii] = buffer[ii];
		//	ii = ii+1;
		//end
		/*
		proc_mem[0] = 8'h30;
		proc_mem[1] = 8'hf4;
		proc_mem[2] = 8'h00;
		proc_mem[3] = 8'h01;
		proc_mem[4] = 8'h00;
		proc_mem[5] = 8'h00;
		proc_mem[6] = 8'h00;
		proc_mem[7] = 8'h00;
		proc_mem[8] = 8'h00;
		proc_mem[9] = 8'h00;
		proc_mem[10] = 8'h00;
		proc_mem[11] = 8'h00;
		proc_mem[12] = 8'h00;
		proc_mem[13] = 8'h00;
		proc_mem[14] = 8'h00;
		*/
		
		
		
proc_mem[0] = 8'h30
;
proc_mem[1] = 8'hf4
;
proc_mem[2] = 8'h00
;
proc_mem[3] = 8'h01
;
proc_mem[4] = 8'h00
;
proc_mem[5] = 8'h00
;
proc_mem[6] = 8'h00
;
proc_mem[7] = 8'h00
;
proc_mem[8] = 8'h00
;
proc_mem[9] = 8'h00
;
proc_mem[10] = 8'h30
;
proc_mem[11] = 8'hf5
;
proc_mem[12] = 8'h00
;
proc_mem[13] = 8'h01
;
proc_mem[14] = 8'h00
;
proc_mem[15] = 8'h00
;
proc_mem[16] = 8'h00
;
proc_mem[17] = 8'h00
;
proc_mem[18] = 8'h00
;
proc_mem[19] = 8'h00
;
proc_mem[20] = 8'h80
;
proc_mem[21] = 8'h40
;
proc_mem[22] = 8'h00
;
proc_mem[23] = 8'h00
;
proc_mem[24] = 8'h00
;
proc_mem[25] = 8'h00
;
proc_mem[26] = 8'h00
;
proc_mem[27] = 8'h00
;
proc_mem[28] = 8'h00
;
proc_mem[29] = 8'h00
;
proc_mem[30] = 8'h00
;
proc_mem[31] = 8'h00
;
proc_mem[32] = 8'h0d
;
proc_mem[33] = 8'h00
;
proc_mem[34] = 8'h00
;
proc_mem[35] = 8'h00
;
proc_mem[36] = 8'h00
;
proc_mem[37] = 8'h00
;
proc_mem[38] = 8'h00
;
proc_mem[39] = 8'h00
;
proc_mem[40] = 8'hc0
;
proc_mem[41] = 8'h00
;
proc_mem[42] = 8'h00
;
proc_mem[43] = 8'h00
;
proc_mem[44] = 8'h00
;
proc_mem[45] = 8'h00
;
proc_mem[46] = 8'h00
;
proc_mem[47] = 8'h00
;
proc_mem[48] = 8'h00
;
proc_mem[49] = 8'h0b
;
proc_mem[50] = 8'h00
;
proc_mem[51] = 8'h00
;
proc_mem[52] = 8'h00
;
proc_mem[53] = 8'h00
;
proc_mem[54] = 8'h00
;
proc_mem[55] = 8'h00
;
proc_mem[56] = 8'h00
;
proc_mem[57] = 8'ha0
;
proc_mem[58] = 8'h00
;
proc_mem[59] = 8'h00
;
proc_mem[60] = 8'h00
;
proc_mem[61] = 8'h00
;
proc_mem[62] = 8'h00
;
proc_mem[63] = 8'h00
;
proc_mem[64] = 8'ha0
;
proc_mem[65] = 8'h5f
;
proc_mem[66] = 8'h20
;
proc_mem[67] = 8'h45
;
proc_mem[68] = 8'h30
;
proc_mem[69] = 8'hf0
;
proc_mem[70] = 8'h04
;
proc_mem[71] = 8'h00
;
proc_mem[72] = 8'h00
;
proc_mem[73] = 8'h00
;
proc_mem[74] = 8'h00
;
proc_mem[75] = 8'h00
;
proc_mem[76] = 8'h00
;
proc_mem[77] = 8'h00
;
proc_mem[78] = 8'ha0
;
proc_mem[79] = 8'h0f
;
proc_mem[80] = 8'h30
;
proc_mem[81] = 8'hf2
;
proc_mem[82] = 8'h20
;
proc_mem[83] = 8'h00
;
proc_mem[84] = 8'h00
;
proc_mem[85] = 8'h00
;
proc_mem[86] = 8'h00
;
proc_mem[87] = 8'h00
;
proc_mem[88] = 8'h00
;
proc_mem[89] = 8'h00
;
proc_mem[90] = 8'ha0
;
proc_mem[91] = 8'h2f
;
proc_mem[92] = 8'h80
;
proc_mem[93] = 8'h6a
;
proc_mem[94] = 8'h00
;
proc_mem[95] = 8'h00
;
proc_mem[96] = 8'h00
;
proc_mem[97] = 8'h00
;
proc_mem[98] = 8'h00
;
proc_mem[99] = 8'h00
;
proc_mem[100] = 8'h00
;
proc_mem[101] = 8'h20
;
proc_mem[102] = 8'h54
;
proc_mem[103] = 8'hb0
;
proc_mem[104] = 8'h5f
;
proc_mem[105] = 8'h90
;
proc_mem[106] = 8'ha0
;
proc_mem[107] = 8'h5f
;
proc_mem[108] = 8'h20
;
proc_mem[109] = 8'h45
;
proc_mem[110] = 8'h50
;
proc_mem[111] = 8'h15
;
proc_mem[112] = 8'h08
;
proc_mem[113] = 8'h00
;
proc_mem[114] = 8'h00
;
proc_mem[115] = 8'h00
;
proc_mem[116] = 8'h00
;
proc_mem[117] = 8'h00
;
proc_mem[118] = 8'h00
;
proc_mem[119] = 8'h00
;
proc_mem[120] = 8'h50
;
proc_mem[121] = 8'h25
;
proc_mem[122] = 8'h0c
;
proc_mem[123] = 8'h00
;
proc_mem[124] = 8'h00
;
proc_mem[125] = 8'h00
;
proc_mem[126] = 8'h00
;
proc_mem[127] = 8'h00
;
proc_mem[128] = 8'h00
;
proc_mem[129] = 8'h00
;
proc_mem[130] = 8'h63
;
proc_mem[131] = 8'h00
;
proc_mem[132] = 8'h62
;
proc_mem[133] = 8'h22
;
proc_mem[134] = 8'h73
;
proc_mem[135] = 8'hbc
;
proc_mem[136] = 8'h00
;
proc_mem[137] = 8'h00
;
proc_mem[138] = 8'h00
;
proc_mem[139] = 8'h00
;
proc_mem[140] = 8'h00
;
proc_mem[141] = 8'h00
;
proc_mem[142] = 8'h00
;
proc_mem[143] = 8'h50
;
proc_mem[144] = 8'h61
;
proc_mem[145] = 8'h00
;
proc_mem[146] = 8'h00
;
proc_mem[147] = 8'h00
;
proc_mem[148] = 8'h00
;
proc_mem[149] = 8'h00
;
proc_mem[150] = 8'h00
;
proc_mem[151] = 8'h00
;
proc_mem[152] = 8'h00
;
proc_mem[153] = 8'h60
;
proc_mem[154] = 8'h60
;
proc_mem[155] = 8'h30
;
proc_mem[156] = 8'hf3
;
proc_mem[157] = 8'h04
;
proc_mem[158] = 8'h00
;
proc_mem[159] = 8'h00
;
proc_mem[160] = 8'h00
;
proc_mem[161] = 8'h00
;
proc_mem[162] = 8'h00
;
proc_mem[163] = 8'h00
;
proc_mem[164] = 8'h00
;
proc_mem[165] = 8'h60
;
proc_mem[166] = 8'h31
;
proc_mem[167] = 8'h30
;
proc_mem[168] = 8'hf3
;
proc_mem[169] = 8'hff
;
proc_mem[170] = 8'hff
;
proc_mem[171] = 8'hff
;
proc_mem[172] = 8'hff
;
proc_mem[173] = 8'hff
;
proc_mem[174] = 8'hff
;
proc_mem[175] = 8'hff
;
proc_mem[176] = 8'hff
;
proc_mem[177] = 8'h60
;
proc_mem[178] = 8'h32
;
proc_mem[179] = 8'h74
;
proc_mem[180] = 8'h8f
;
proc_mem[181] = 8'h00
;
proc_mem[182] = 8'h00
;
proc_mem[183] = 8'h00
;
proc_mem[184] = 8'h00
;
proc_mem[185] = 8'h00
;
proc_mem[186] = 8'h00
;
proc_mem[187] = 8'h00
;
proc_mem[188] = 8'h20
;
proc_mem[189] = 8'h54
;
proc_mem[190] = 8'hb0
;
proc_mem[191] = 8'h5f
;
proc_mem[192] = 8'h90
;
proc_mem[193] = 8'h90
;
proc_mem[194] = 8'h00;
proc_mem[195] = 8'h00;
proc_mem[196] = 8'h00;
proc_mem[197] = 8'h00;
proc_mem[198] = 8'h00;
proc_mem[199] = 8'h00;
proc_mem[200] = 8'h00;
proc_mem[201] = 8'h00;
proc_mem[202] = 8'h00;
proc_mem[203] = 8'h00;
proc_mem[204] = 8'h00;
proc_mem[205] = 8'h00;
proc_mem[206] = 8'h00;
proc_mem[207] = 8'h00;
proc_mem[208] = 8'h00;
proc_mem[209] = 8'h00;
proc_mem[210] = 8'h00;
proc_mem[211] = 8'h00;
proc_mem[212] = 8'h00;
proc_mem[213] = 8'h00;
proc_mem[214] = 8'h00;
proc_mem[215] = 8'h00;
proc_mem[216] = 8'h00;
proc_mem[217] = 8'h00;
proc_mem[218] = 8'h00;
proc_mem[219] = 8'h00;
proc_mem[220] = 8'h00;
proc_mem[221] = 8'h00;
proc_mem[222] = 8'h00;
proc_mem[223] = 8'h00;
proc_mem[224] = 8'h00;
proc_mem[225] = 8'h00;
proc_mem[226] = 8'h00;
proc_mem[227] = 8'h00;
proc_mem[228] = 8'h00;
proc_mem[229] = 8'h00;
proc_mem[230] = 8'h00;
proc_mem[231] = 8'h00;
proc_mem[232] = 8'h00;
proc_mem[233] = 8'h00;
proc_mem[234] = 8'h00;
proc_mem[235] = 8'h00;
proc_mem[236] = 8'h00;
proc_mem[237] = 8'h00;
proc_mem[238] = 8'h00;
proc_mem[239] = 8'h00;
proc_mem[240] = 8'h00;
proc_mem[241] = 8'h00;
proc_mem[242] = 8'h00;
proc_mem[243] = 8'h00;
proc_mem[244] = 8'h00;
proc_mem[245] = 8'h00;
proc_mem[246] = 8'h00;
proc_mem[247] = 8'h00;
proc_mem[248] = 8'h00;
proc_mem[249] = 8'h00;
proc_mem[250] = 8'h00;
proc_mem[251] = 8'h00;
proc_mem[252] = 8'h00;
proc_mem[253] = 8'h00;
proc_mem[254] = 8'h00;
proc_mem[255] = 8'h00;
proc_mem[256] = 8'h00;
proc_mem[257] = 8'h00;
proc_mem[258] = 8'h00;
proc_mem[259] = 8'h00;
proc_mem[260] = 8'h00;
proc_mem[261] = 8'h00;
proc_mem[262] = 8'h00;
proc_mem[263] = 8'h00;
proc_mem[264] = 8'h00;
proc_mem[265] = 8'h00;
proc_mem[266] = 8'h00;
proc_mem[267] = 8'h00;
proc_mem[268] = 8'h00;
proc_mem[269] = 8'h00;
proc_mem[270] = 8'h00;
proc_mem[271] = 8'h00;
proc_mem[272] = 8'h00;
proc_mem[273] = 8'h00;
proc_mem[274] = 8'h00;
proc_mem[275] = 8'h00;
proc_mem[276] = 8'h00;
proc_mem[277] = 8'h00;
proc_mem[278] = 8'h00;
proc_mem[279] = 8'h00;
proc_mem[280] = 8'h00;
proc_mem[281] = 8'h00;
proc_mem[282] = 8'h00;
proc_mem[283] = 8'h00;
proc_mem[284] = 8'h00;
proc_mem[285] = 8'h00;
proc_mem[286] = 8'h00;
proc_mem[287] = 8'h00;
proc_mem[288] = 8'h00;
proc_mem[289] = 8'h00;
proc_mem[290] = 8'h00;
proc_mem[291] = 8'h00;
proc_mem[292] = 8'h00;
proc_mem[293] = 8'h00;
proc_mem[294] = 8'h00;
proc_mem[295] = 8'h00;
proc_mem[296] = 8'h00;
proc_mem[297] = 8'h00;
proc_mem[298] = 8'h00;
proc_mem[299] = 8'h00;
proc_mem[300] = 8'h00;
proc_mem[301] = 8'h00;
proc_mem[302] = 8'h00;
proc_mem[303] = 8'h00;
proc_mem[304] = 8'h00;
proc_mem[305] = 8'h00;
proc_mem[306] = 8'h00;
proc_mem[307] = 8'h00;
proc_mem[308] = 8'h00;
proc_mem[309] = 8'h00;
proc_mem[310] = 8'h00;
proc_mem[311] = 8'h00;
proc_mem[312] = 8'h00;
proc_mem[313] = 8'h00;
proc_mem[314] = 8'h00;
proc_mem[315] = 8'h00;
proc_mem[316] = 8'h00;
proc_mem[317] = 8'h00;
proc_mem[318] = 8'h00;
proc_mem[319] = 8'h00;
proc_mem[320] = 8'h00;
proc_mem[321] = 8'h00;
proc_mem[322] = 8'h00;
proc_mem[323] = 8'h00;
proc_mem[324] = 8'h00;
proc_mem[325] = 8'h00;
proc_mem[326] = 8'h00;
proc_mem[327] = 8'h00;
proc_mem[328] = 8'h00;
proc_mem[329] = 8'h00;
proc_mem[330] = 8'h00;
proc_mem[331] = 8'h00;
proc_mem[332] = 8'h00;
proc_mem[333] = 8'h00;
proc_mem[334] = 8'h00;
proc_mem[335] = 8'h00;
proc_mem[336] = 8'h00;
proc_mem[337] = 8'h00;
proc_mem[338] = 8'h00;
proc_mem[339] = 8'h00;
proc_mem[340] = 8'h00;
proc_mem[341] = 8'h00;
proc_mem[342] = 8'h00;
proc_mem[343] = 8'h00;
proc_mem[344] = 8'h00;
proc_mem[345] = 8'h00;
proc_mem[346] = 8'h00;
proc_mem[347] = 8'h00;
proc_mem[348] = 8'h00;
proc_mem[349] = 8'h00;
proc_mem[350] = 8'h00;
proc_mem[351] = 8'h00;
proc_mem[352] = 8'h00;
proc_mem[353] = 8'h00;
proc_mem[354] = 8'h00;
proc_mem[355] = 8'h00;
proc_mem[356] = 8'h00;
proc_mem[357] = 8'h00;
proc_mem[358] = 8'h00;
proc_mem[359] = 8'h00;
proc_mem[360] = 8'h00;
proc_mem[361] = 8'h00;
proc_mem[362] = 8'h00;
proc_mem[363] = 8'h00;
proc_mem[364] = 8'h00;
proc_mem[365] = 8'h00;
proc_mem[366] = 8'h00;
proc_mem[367] = 8'h00;
proc_mem[368] = 8'h00;
proc_mem[369] = 8'h00;
proc_mem[370] = 8'h00;
proc_mem[371] = 8'h00;
proc_mem[372] = 8'h00;
proc_mem[373] = 8'h00;
proc_mem[374] = 8'h00;
proc_mem[375] = 8'h00;
proc_mem[376] = 8'h00;
proc_mem[377] = 8'h00;
proc_mem[378] = 8'h00;
proc_mem[379] = 8'h00;
proc_mem[380] = 8'h00;
proc_mem[381] = 8'h00;
proc_mem[382] = 8'h00;
proc_mem[383] = 8'h00;
proc_mem[384] = 8'h00;
proc_mem[385] = 8'h00;
proc_mem[386] = 8'h00;
proc_mem[387] = 8'h00;
proc_mem[388] = 8'h00;
proc_mem[389] = 8'h00;
proc_mem[390] = 8'h00;
proc_mem[391] = 8'h00;
proc_mem[392] = 8'h00;
proc_mem[393] = 8'h00;
proc_mem[394] = 8'h00;
proc_mem[395] = 8'h00;
proc_mem[396] = 8'h00;
proc_mem[397] = 8'h00;
proc_mem[398] = 8'h00;
proc_mem[399] = 8'h00;
proc_mem[400] = 8'h00;
proc_mem[401] = 8'h00;
proc_mem[402] = 8'h00;
proc_mem[403] = 8'h00;
proc_mem[404] = 8'h00;
proc_mem[405] = 8'h00;
proc_mem[406] = 8'h00;
proc_mem[407] = 8'h00;
proc_mem[408] = 8'h00;
proc_mem[409] = 8'h00;
proc_mem[410] = 8'h00;
proc_mem[411] = 8'h00;
proc_mem[412] = 8'h00;
proc_mem[413] = 8'h00;
proc_mem[414] = 8'h00;
proc_mem[415] = 8'h00;
proc_mem[416] = 8'h00;
proc_mem[417] = 8'h00;
proc_mem[418] = 8'h00;
proc_mem[419] = 8'h00;
proc_mem[420] = 8'h00;
proc_mem[421] = 8'h00;
proc_mem[422] = 8'h00;
proc_mem[423] = 8'h00;
proc_mem[424] = 8'h00;
proc_mem[425] = 8'h00;
proc_mem[426] = 8'h00;
proc_mem[427] = 8'h00;
proc_mem[428] = 8'h00;
proc_mem[429] = 8'h00;
proc_mem[430] = 8'h00;
proc_mem[431] = 8'h00;
proc_mem[432] = 8'h00;
proc_mem[433] = 8'h00;
proc_mem[434] = 8'h00;
proc_mem[435] = 8'h00;
proc_mem[436] = 8'h00;
proc_mem[437] = 8'h00;
proc_mem[438] = 8'h00;
proc_mem[439] = 8'h00;
proc_mem[440] = 8'h00;
proc_mem[441] = 8'h00;
proc_mem[442] = 8'h00;
proc_mem[443] = 8'h00;
proc_mem[444] = 8'h00;
proc_mem[445] = 8'h00;
proc_mem[446] = 8'h00;
proc_mem[447] = 8'h00;
proc_mem[448] = 8'h00;
proc_mem[449] = 8'h00;
proc_mem[450] = 8'h00;
proc_mem[451] = 8'h00;
proc_mem[452] = 8'h00;
proc_mem[453] = 8'h00;
proc_mem[454] = 8'h00;
proc_mem[455] = 8'h00;
proc_mem[456] = 8'h00;
proc_mem[457] = 8'h00;
proc_mem[458] = 8'h00;
proc_mem[459] = 8'h00;
proc_mem[460] = 8'h00;
proc_mem[461] = 8'h00;
proc_mem[462] = 8'h00;
proc_mem[463] = 8'h00;
proc_mem[464] = 8'h00;
proc_mem[465] = 8'h00;
proc_mem[466] = 8'h00;
proc_mem[467] = 8'h00;
proc_mem[468] = 8'h00;
proc_mem[469] = 8'h00;
proc_mem[470] = 8'h00;
proc_mem[471] = 8'h00;
proc_mem[472] = 8'h00;
proc_mem[473] = 8'h00;
proc_mem[474] = 8'h00;
proc_mem[475] = 8'h00;
proc_mem[476] = 8'h00;
proc_mem[477] = 8'h00;
proc_mem[478] = 8'h00;
proc_mem[479] = 8'h00;
proc_mem[480] = 8'h00;
proc_mem[481] = 8'h00;
proc_mem[482] = 8'h00;
proc_mem[483] = 8'h00;
proc_mem[484] = 8'h00;
proc_mem[485] = 8'h00;
proc_mem[486] = 8'h00;
proc_mem[487] = 8'h00;
proc_mem[488] = 8'h00;
proc_mem[489] = 8'h00;
proc_mem[490] = 8'h00;
proc_mem[491] = 8'h00;
proc_mem[492] = 8'h00;
proc_mem[493] = 8'h00;
proc_mem[494] = 8'h00;
proc_mem[495] = 8'h00;
proc_mem[496] = 8'h00;
proc_mem[497] = 8'h00;
proc_mem[498] = 8'h00;
proc_mem[499] = 8'h00;
proc_mem[500] = 8'h00;
proc_mem[501] = 8'h00;
proc_mem[502] = 8'h00;
proc_mem[503] = 8'h00;
proc_mem[504] = 8'h00;
proc_mem[505] = 8'h00;
proc_mem[506] = 8'h00;
proc_mem[507] = 8'h00;
proc_mem[508] = 8'h00;
proc_mem[509] = 8'h00;
proc_mem[510] = 8'h00;
proc_mem[511] = 8'h00;
proc_mem[512] = 8'h00;
proc_mem[513] = 8'h00;
proc_mem[514] = 8'h00;
proc_mem[515] = 8'h00;
proc_mem[516] = 8'h00;
proc_mem[517] = 8'h00;
proc_mem[518] = 8'h00;
proc_mem[519] = 8'h00;
proc_mem[520] = 8'h00;
proc_mem[521] = 8'h00;
proc_mem[522] = 8'h00;
proc_mem[523] = 8'h00;
proc_mem[524] = 8'h00;
proc_mem[525] = 8'h00;
proc_mem[526] = 8'h00;
proc_mem[527] = 8'h00;
proc_mem[528] = 8'h00;
proc_mem[529] = 8'h00;
proc_mem[530] = 8'h00;
proc_mem[531] = 8'h00;
proc_mem[532] = 8'h00;
proc_mem[533] = 8'h00;
proc_mem[534] = 8'h00;
proc_mem[535] = 8'h00;
proc_mem[536] = 8'h00;
proc_mem[537] = 8'h00;
proc_mem[538] = 8'h00;
proc_mem[539] = 8'h00;
proc_mem[540] = 8'h00;
proc_mem[541] = 8'h00;
proc_mem[542] = 8'h00;
proc_mem[543] = 8'h00;
proc_mem[544] = 8'h00;
proc_mem[545] = 8'h00;
proc_mem[546] = 8'h00;
proc_mem[547] = 8'h00;
proc_mem[548] = 8'h00;
proc_mem[549] = 8'h00;
proc_mem[550] = 8'h00;
proc_mem[551] = 8'h00;
proc_mem[552] = 8'h00;
proc_mem[553] = 8'h00;
proc_mem[554] = 8'h00;
proc_mem[555] = 8'h00;
proc_mem[556] = 8'h00;
proc_mem[557] = 8'h00;
proc_mem[558] = 8'h00;
proc_mem[559] = 8'h00;
proc_mem[560] = 8'h00;
proc_mem[561] = 8'h00;
proc_mem[562] = 8'h00;
proc_mem[563] = 8'h00;
proc_mem[564] = 8'h00;
proc_mem[565] = 8'h00;
proc_mem[566] = 8'h00;
proc_mem[567] = 8'h00;
proc_mem[568] = 8'h00;
proc_mem[569] = 8'h00;
proc_mem[570] = 8'h00;
proc_mem[571] = 8'h00;
proc_mem[572] = 8'h00;
proc_mem[573] = 8'h00;
proc_mem[574] = 8'h00;
proc_mem[575] = 8'h00;
proc_mem[576] = 8'h00;
proc_mem[577] = 8'h00;
proc_mem[578] = 8'h00;
proc_mem[579] = 8'h00;
proc_mem[580] = 8'h00;
proc_mem[581] = 8'h00;
proc_mem[582] = 8'h00;
proc_mem[583] = 8'h00;
proc_mem[584] = 8'h00;
proc_mem[585] = 8'h00;
proc_mem[586] = 8'h00;
proc_mem[587] = 8'h00;
proc_mem[588] = 8'h00;
proc_mem[589] = 8'h00;
proc_mem[590] = 8'h00;
proc_mem[591] = 8'h00;
proc_mem[592] = 8'h00;
proc_mem[593] = 8'h00;
proc_mem[594] = 8'h00;
proc_mem[595] = 8'h00;
proc_mem[596] = 8'h00;
proc_mem[597] = 8'h00;
proc_mem[598] = 8'h00;
proc_mem[599] = 8'h00;
proc_mem[600] = 8'h00;
proc_mem[601] = 8'h00;
proc_mem[602] = 8'h00;
proc_mem[603] = 8'h00;
proc_mem[604] = 8'h00;
proc_mem[605] = 8'h00;
proc_mem[606] = 8'h00;
proc_mem[607] = 8'h00;
proc_mem[608] = 8'h00;
proc_mem[609] = 8'h00;
proc_mem[610] = 8'h00;
proc_mem[611] = 8'h00;
proc_mem[612] = 8'h00;
proc_mem[613] = 8'h00;
proc_mem[614] = 8'h00;
proc_mem[615] = 8'h00;
proc_mem[616] = 8'h00;
proc_mem[617] = 8'h00;
proc_mem[618] = 8'h00;
proc_mem[619] = 8'h00;
proc_mem[620] = 8'h00;
proc_mem[621] = 8'h00;
proc_mem[622] = 8'h00;
proc_mem[623] = 8'h00;
proc_mem[624] = 8'h00;
proc_mem[625] = 8'h00;
proc_mem[626] = 8'h00;
proc_mem[627] = 8'h00;
proc_mem[628] = 8'h00;
proc_mem[629] = 8'h00;
proc_mem[630] = 8'h00;
proc_mem[631] = 8'h00;
proc_mem[632] = 8'h00;
proc_mem[633] = 8'h00;
proc_mem[634] = 8'h00;
proc_mem[635] = 8'h00;
proc_mem[636] = 8'h00;
proc_mem[637] = 8'h00;
proc_mem[638] = 8'h00;
proc_mem[639] = 8'h00;
proc_mem[640] = 8'h00;
proc_mem[641] = 8'h00;
proc_mem[642] = 8'h00;
proc_mem[643] = 8'h00;
proc_mem[644] = 8'h00;
proc_mem[645] = 8'h00;
proc_mem[646] = 8'h00;
proc_mem[647] = 8'h00;
proc_mem[648] = 8'h00;
proc_mem[649] = 8'h00;
proc_mem[650] = 8'h00;
proc_mem[651] = 8'h00;
proc_mem[652] = 8'h00;
proc_mem[653] = 8'h00;
proc_mem[654] = 8'h00;
proc_mem[655] = 8'h00;
proc_mem[656] = 8'h00;
proc_mem[657] = 8'h00;
proc_mem[658] = 8'h00;
proc_mem[659] = 8'h00;
proc_mem[660] = 8'h00;
proc_mem[661] = 8'h00;
proc_mem[662] = 8'h00;
proc_mem[663] = 8'h00;
proc_mem[664] = 8'h00;
proc_mem[665] = 8'h00;
proc_mem[666] = 8'h00;
proc_mem[667] = 8'h00;
proc_mem[668] = 8'h00;
proc_mem[669] = 8'h00;
proc_mem[670] = 8'h00;
proc_mem[671] = 8'h00;
proc_mem[672] = 8'h00;
proc_mem[673] = 8'h00;
proc_mem[674] = 8'h00;
proc_mem[675] = 8'h00;
proc_mem[676] = 8'h00;
proc_mem[677] = 8'h00;
proc_mem[678] = 8'h00;
proc_mem[679] = 8'h00;
proc_mem[680] = 8'h00;
proc_mem[681] = 8'h00;
proc_mem[682] = 8'h00;
proc_mem[683] = 8'h00;
proc_mem[684] = 8'h00;
proc_mem[685] = 8'h00;
proc_mem[686] = 8'h00;
proc_mem[687] = 8'h00;
proc_mem[688] = 8'h00;
proc_mem[689] = 8'h00;
proc_mem[690] = 8'h00;
proc_mem[691] = 8'h00;
proc_mem[692] = 8'h00;
proc_mem[693] = 8'h00;
proc_mem[694] = 8'h00;
proc_mem[695] = 8'h00;
proc_mem[696] = 8'h00;
proc_mem[697] = 8'h00;
proc_mem[698] = 8'h00;
proc_mem[699] = 8'h00;
proc_mem[700] = 8'h00;
proc_mem[701] = 8'h00;
proc_mem[702] = 8'h00;
proc_mem[703] = 8'h00;
proc_mem[704] = 8'h00;
proc_mem[705] = 8'h00;
proc_mem[706] = 8'h00;
proc_mem[707] = 8'h00;
proc_mem[708] = 8'h00;
proc_mem[709] = 8'h00;
proc_mem[710] = 8'h00;
proc_mem[711] = 8'h00;
proc_mem[712] = 8'h00;
proc_mem[713] = 8'h00;
proc_mem[714] = 8'h00;
proc_mem[715] = 8'h00;
proc_mem[716] = 8'h00;
proc_mem[717] = 8'h00;
proc_mem[718] = 8'h00;
proc_mem[719] = 8'h00;
proc_mem[720] = 8'h00;
proc_mem[721] = 8'h00;
proc_mem[722] = 8'h00;
proc_mem[723] = 8'h00;
proc_mem[724] = 8'h00;
proc_mem[725] = 8'h00;
proc_mem[726] = 8'h00;
proc_mem[727] = 8'h00;
proc_mem[728] = 8'h00;
proc_mem[729] = 8'h00;
proc_mem[730] = 8'h00;
proc_mem[731] = 8'h00;
proc_mem[732] = 8'h00;
proc_mem[733] = 8'h00;
proc_mem[734] = 8'h00;
proc_mem[735] = 8'h00;
proc_mem[736] = 8'h00;
proc_mem[737] = 8'h00;
proc_mem[738] = 8'h00;
proc_mem[739] = 8'h00;
proc_mem[740] = 8'h00;
proc_mem[741] = 8'h00;
proc_mem[742] = 8'h00;
proc_mem[743] = 8'h00;
proc_mem[744] = 8'h00;
proc_mem[745] = 8'h00;
proc_mem[746] = 8'h00;
proc_mem[747] = 8'h00;
proc_mem[748] = 8'h00;
proc_mem[749] = 8'h00;
proc_mem[750] = 8'h00;
proc_mem[751] = 8'h00;
proc_mem[752] = 8'h00;
proc_mem[753] = 8'h00;
proc_mem[754] = 8'h00;
proc_mem[755] = 8'h00;
proc_mem[756] = 8'h00;
proc_mem[757] = 8'h00;
proc_mem[758] = 8'h00;
proc_mem[759] = 8'h00;
proc_mem[760] = 8'h00;
proc_mem[761] = 8'h00;
proc_mem[762] = 8'h00;
proc_mem[763] = 8'h00;
proc_mem[764] = 8'h00;
proc_mem[765] = 8'h00;
proc_mem[766] = 8'h00;
proc_mem[767] = 8'h00;
proc_mem[768] = 8'h00;
proc_mem[769] = 8'h00;
proc_mem[770] = 8'h00;
proc_mem[771] = 8'h00;
proc_mem[772] = 8'h00;
proc_mem[773] = 8'h00;
proc_mem[774] = 8'h00;
proc_mem[775] = 8'h00;
proc_mem[776] = 8'h00;
proc_mem[777] = 8'h00;
proc_mem[778] = 8'h00;
proc_mem[779] = 8'h00;
proc_mem[780] = 8'h00;
proc_mem[781] = 8'h00;
proc_mem[782] = 8'h00;
proc_mem[783] = 8'h00;
proc_mem[784] = 8'h00;
proc_mem[785] = 8'h00;
proc_mem[786] = 8'h00;
proc_mem[787] = 8'h00;
proc_mem[788] = 8'h00;
proc_mem[789] = 8'h00;
proc_mem[790] = 8'h00;
proc_mem[791] = 8'h00;
proc_mem[792] = 8'h00;
proc_mem[793] = 8'h00;
proc_mem[794] = 8'h00;
proc_mem[795] = 8'h00;
proc_mem[796] = 8'h00;
proc_mem[797] = 8'h00;
proc_mem[798] = 8'h00;
proc_mem[799] = 8'h00;
proc_mem[800] = 8'h00;
proc_mem[801] = 8'h00;
proc_mem[802] = 8'h00;
proc_mem[803] = 8'h00;
proc_mem[804] = 8'h00;
proc_mem[805] = 8'h00;
proc_mem[806] = 8'h00;
proc_mem[807] = 8'h00;
proc_mem[808] = 8'h00;
proc_mem[809] = 8'h00;
proc_mem[810] = 8'h00;
proc_mem[811] = 8'h00;
proc_mem[812] = 8'h00;
proc_mem[813] = 8'h00;
proc_mem[814] = 8'h00;
proc_mem[815] = 8'h00;
proc_mem[816] = 8'h00;
proc_mem[817] = 8'h00;
proc_mem[818] = 8'h00;
proc_mem[819] = 8'h00;
proc_mem[820] = 8'h00;
proc_mem[821] = 8'h00;
proc_mem[822] = 8'h00;
proc_mem[823] = 8'h00;
proc_mem[824] = 8'h00;
proc_mem[825] = 8'h00;
proc_mem[826] = 8'h00;
proc_mem[827] = 8'h00;
proc_mem[828] = 8'h00;
proc_mem[829] = 8'h00;
proc_mem[830] = 8'h00;
proc_mem[831] = 8'h00;
proc_mem[832] = 8'h00;
proc_mem[833] = 8'h00;
proc_mem[834] = 8'h00;
proc_mem[835] = 8'h00;
proc_mem[836] = 8'h00;
proc_mem[837] = 8'h00;
proc_mem[838] = 8'h00;
proc_mem[839] = 8'h00;
proc_mem[840] = 8'h00;
proc_mem[841] = 8'h00;
proc_mem[842] = 8'h00;
proc_mem[843] = 8'h00;
proc_mem[844] = 8'h00;
proc_mem[845] = 8'h00;
proc_mem[846] = 8'h00;
proc_mem[847] = 8'h00;
proc_mem[848] = 8'h00;
proc_mem[849] = 8'h00;
proc_mem[850] = 8'h00;
proc_mem[851] = 8'h00;
proc_mem[852] = 8'h00;
proc_mem[853] = 8'h00;
proc_mem[854] = 8'h00;
proc_mem[855] = 8'h00;
proc_mem[856] = 8'h00;
proc_mem[857] = 8'h00;
proc_mem[858] = 8'h00;
proc_mem[859] = 8'h00;
proc_mem[860] = 8'h00;
proc_mem[861] = 8'h00;
proc_mem[862] = 8'h00;
proc_mem[863] = 8'h00;
proc_mem[864] = 8'h00;
proc_mem[865] = 8'h00;
proc_mem[866] = 8'h00;
proc_mem[867] = 8'h00;
proc_mem[868] = 8'h00;
proc_mem[869] = 8'h00;
proc_mem[870] = 8'h00;
proc_mem[871] = 8'h00;
proc_mem[872] = 8'h00;
proc_mem[873] = 8'h00;
proc_mem[874] = 8'h00;
proc_mem[875] = 8'h00;
proc_mem[876] = 8'h00;
proc_mem[877] = 8'h00;
proc_mem[878] = 8'h00;
proc_mem[879] = 8'h00;
proc_mem[880] = 8'h00;
proc_mem[881] = 8'h00;
proc_mem[882] = 8'h00;
proc_mem[883] = 8'h00;
proc_mem[884] = 8'h00;
proc_mem[885] = 8'h00;
proc_mem[886] = 8'h00;
proc_mem[887] = 8'h00;
proc_mem[888] = 8'h00;
proc_mem[889] = 8'h00;
proc_mem[890] = 8'h00;
proc_mem[891] = 8'h00;
proc_mem[892] = 8'h00;
proc_mem[893] = 8'h00;
proc_mem[894] = 8'h00;
proc_mem[895] = 8'h00;
proc_mem[896] = 8'h00;
proc_mem[897] = 8'h00;
proc_mem[898] = 8'h00;
proc_mem[899] = 8'h00;
proc_mem[900] = 8'h00;
proc_mem[901] = 8'h00;
proc_mem[902] = 8'h00;
proc_mem[903] = 8'h00;
proc_mem[904] = 8'h00;
proc_mem[905] = 8'h00;
proc_mem[906] = 8'h00;
proc_mem[907] = 8'h00;
proc_mem[908] = 8'h00;
proc_mem[909] = 8'h00;
proc_mem[910] = 8'h00;
proc_mem[911] = 8'h00;
proc_mem[912] = 8'h00;
proc_mem[913] = 8'h00;
proc_mem[914] = 8'h00;
proc_mem[915] = 8'h00;
proc_mem[916] = 8'h00;
proc_mem[917] = 8'h00;
proc_mem[918] = 8'h00;
proc_mem[919] = 8'h00;
proc_mem[920] = 8'h00;
proc_mem[921] = 8'h00;
proc_mem[922] = 8'h00;
proc_mem[923] = 8'h00;
proc_mem[924] = 8'h00;
proc_mem[925] = 8'h00;
proc_mem[926] = 8'h00;
proc_mem[927] = 8'h00;
proc_mem[928] = 8'h00;
proc_mem[929] = 8'h00;
proc_mem[930] = 8'h00;
proc_mem[931] = 8'h00;
proc_mem[932] = 8'h00;
proc_mem[933] = 8'h00;
proc_mem[934] = 8'h00;
proc_mem[935] = 8'h00;
proc_mem[936] = 8'h00;
proc_mem[937] = 8'h00;
proc_mem[938] = 8'h00;
proc_mem[939] = 8'h00;
proc_mem[940] = 8'h00;
proc_mem[941] = 8'h00;
proc_mem[942] = 8'h00;
proc_mem[943] = 8'h00;
proc_mem[944] = 8'h00;
proc_mem[945] = 8'h00;
proc_mem[946] = 8'h00;
proc_mem[947] = 8'h00;
proc_mem[948] = 8'h00;
proc_mem[949] = 8'h00;
proc_mem[950] = 8'h00;
proc_mem[951] = 8'h00;
proc_mem[952] = 8'h00;
proc_mem[953] = 8'h00;
proc_mem[954] = 8'h00;
proc_mem[955] = 8'h00;
proc_mem[956] = 8'h00;
proc_mem[957] = 8'h00;
proc_mem[958] = 8'h00;
proc_mem[959] = 8'h00;
proc_mem[960] = 8'h00;
proc_mem[961] = 8'h00;
proc_mem[962] = 8'h00;
proc_mem[963] = 8'h00;
proc_mem[964] = 8'h00;
proc_mem[965] = 8'h00;
proc_mem[966] = 8'h00;
proc_mem[967] = 8'h00;
proc_mem[968] = 8'h00;
proc_mem[969] = 8'h00;
proc_mem[970] = 8'h00;
proc_mem[971] = 8'h00;
proc_mem[972] = 8'h00;
proc_mem[973] = 8'h00;
proc_mem[974] = 8'h00;
proc_mem[975] = 8'h00;
proc_mem[976] = 8'h00;
proc_mem[977] = 8'h00;
proc_mem[978] = 8'h00;
proc_mem[979] = 8'h00;
proc_mem[980] = 8'h00;
proc_mem[981] = 8'h00;
proc_mem[982] = 8'h00;
proc_mem[983] = 8'h00;
proc_mem[984] = 8'h00;
proc_mem[985] = 8'h00;
proc_mem[986] = 8'h00;
proc_mem[987] = 8'h00;
proc_mem[988] = 8'h00;
proc_mem[989] = 8'h00;
proc_mem[990] = 8'h00;
proc_mem[991] = 8'h00;
proc_mem[992] = 8'h00;
proc_mem[993] = 8'h00;
proc_mem[994] = 8'h00;
proc_mem[995] = 8'h00;
proc_mem[996] = 8'h00;
proc_mem[997] = 8'h00;
proc_mem[998] = 8'h00;
proc_mem[999] = 8'h00;
proc_mem[1000] = 8'h00;
proc_mem[1001] = 8'h00;
proc_mem[1002] = 8'h00;
proc_mem[1003] = 8'h00;
proc_mem[1004] = 8'h00;
proc_mem[1005] = 8'h00;
proc_mem[1006] = 8'h00;
proc_mem[1007] = 8'h00;
proc_mem[1008] = 8'h00;
proc_mem[1009] = 8'h00;
proc_mem[1010] = 8'h00;
proc_mem[1011] = 8'h00;
proc_mem[1012] = 8'h00;
proc_mem[1013] = 8'h00;
proc_mem[1014] = 8'h00;
proc_mem[1015] = 8'h00;
proc_mem[1016] = 8'h00;
proc_mem[1017] = 8'h00;
proc_mem[1018] = 8'h00;
proc_mem[1019] = 8'h00;
proc_mem[1020] = 8'h00;
proc_mem[1021] = 8'h00;
proc_mem[1022] = 8'h00;
proc_mem[1023] = 8'h00;
proc_mem[1024] = 8'h00;
proc_mem[1025] = 8'h00;
proc_mem[1026] = 8'h00;
proc_mem[1027] = 8'h00;
proc_mem[1028] = 8'h00;
proc_mem[1029] = 8'h00;
proc_mem[1030] = 8'h00;
proc_mem[1031] = 8'h00;
proc_mem[1032] = 8'h00;
proc_mem[1033] = 8'h00;
proc_mem[1034] = 8'h00;
proc_mem[1035] = 8'h00;
proc_mem[1036] = 8'h00;
proc_mem[1037] = 8'h00;
proc_mem[1038] = 8'h00;
proc_mem[1039] = 8'h00;
proc_mem[1040] = 8'h00;
proc_mem[1041] = 8'h00;
proc_mem[1042] = 8'h00;
proc_mem[1043] = 8'h00;
proc_mem[1044] = 8'h00;
proc_mem[1045] = 8'h00;
proc_mem[1046] = 8'h00;
proc_mem[1047] = 8'h00;
proc_mem[1048] = 8'h00;
proc_mem[1049] = 8'h00;
proc_mem[1050] = 8'h00;
proc_mem[1051] = 8'h00;
proc_mem[1052] = 8'h00;
proc_mem[1053] = 8'h00;
proc_mem[1054] = 8'h00;
proc_mem[1055] = 8'h00;
proc_mem[1056] = 8'h00;
proc_mem[1057] = 8'h00;
proc_mem[1058] = 8'h00;
proc_mem[1059] = 8'h00;
proc_mem[1060] = 8'h00;
proc_mem[1061] = 8'h00;
proc_mem[1062] = 8'h00;
proc_mem[1063] = 8'h00;
proc_mem[1064] = 8'h00;
proc_mem[1065] = 8'h00;
proc_mem[1066] = 8'h00;
proc_mem[1067] = 8'h00;
proc_mem[1068] = 8'h00;
proc_mem[1069] = 8'h00;
proc_mem[1070] = 8'h00;
proc_mem[1071] = 8'h00;
proc_mem[1072] = 8'h00;
proc_mem[1073] = 8'h00;
proc_mem[1074] = 8'h00;
proc_mem[1075] = 8'h00;
proc_mem[1076] = 8'h00;
proc_mem[1077] = 8'h00;
proc_mem[1078] = 8'h00;
proc_mem[1079] = 8'h00;
proc_mem[1080] = 8'h00;
proc_mem[1081] = 8'h00;
proc_mem[1082] = 8'h00;
proc_mem[1083] = 8'h00;
proc_mem[1084] = 8'h00;
proc_mem[1085] = 8'h00;
proc_mem[1086] = 8'h00;
proc_mem[1087] = 8'h00;
proc_mem[1088] = 8'h00;
proc_mem[1089] = 8'h00;
proc_mem[1090] = 8'h00;
proc_mem[1091] = 8'h00;
proc_mem[1092] = 8'h00;
proc_mem[1093] = 8'h00;
proc_mem[1094] = 8'h00;
proc_mem[1095] = 8'h00;
proc_mem[1096] = 8'h00;
proc_mem[1097] = 8'h00;
proc_mem[1098] = 8'h00;
proc_mem[1099] = 8'h00;
proc_mem[1100] = 8'h00;
proc_mem[1101] = 8'h00;
proc_mem[1102] = 8'h00;
proc_mem[1103] = 8'h00;
proc_mem[1104] = 8'h00;
proc_mem[1105] = 8'h00;
proc_mem[1106] = 8'h00;
proc_mem[1107] = 8'h00;
proc_mem[1108] = 8'h00;
proc_mem[1109] = 8'h00;
proc_mem[1110] = 8'h00;
proc_mem[1111] = 8'h00;
proc_mem[1112] = 8'h00;
proc_mem[1113] = 8'h00;
proc_mem[1114] = 8'h00;
proc_mem[1115] = 8'h00;
proc_mem[1116] = 8'h00;
proc_mem[1117] = 8'h00;
proc_mem[1118] = 8'h00;
proc_mem[1119] = 8'h00;
proc_mem[1120] = 8'h00;
proc_mem[1121] = 8'h00;
proc_mem[1122] = 8'h00;
proc_mem[1123] = 8'h00;
proc_mem[1124] = 8'h00;
proc_mem[1125] = 8'h00;
proc_mem[1126] = 8'h00;
proc_mem[1127] = 8'h00;
proc_mem[1128] = 8'h00;
proc_mem[1129] = 8'h00;
proc_mem[1130] = 8'h00;
proc_mem[1131] = 8'h00;
proc_mem[1132] = 8'h00;
proc_mem[1133] = 8'h00;
proc_mem[1134] = 8'h00;
proc_mem[1135] = 8'h00;
proc_mem[1136] = 8'h00;
proc_mem[1137] = 8'h00;
proc_mem[1138] = 8'h00;
proc_mem[1139] = 8'h00;
proc_mem[1140] = 8'h00;
proc_mem[1141] = 8'h00;
proc_mem[1142] = 8'h00;
proc_mem[1143] = 8'h00;
proc_mem[1144] = 8'h00;
proc_mem[1145] = 8'h00;
proc_mem[1146] = 8'h00;
proc_mem[1147] = 8'h00;
proc_mem[1148] = 8'h00;
proc_mem[1149] = 8'h00;
proc_mem[1150] = 8'h00;
proc_mem[1151] = 8'h00;
proc_mem[1152] = 8'h00;
proc_mem[1153] = 8'h00;
proc_mem[1154] = 8'h00;
proc_mem[1155] = 8'h00;
proc_mem[1156] = 8'h00;
proc_mem[1157] = 8'h00;
proc_mem[1158] = 8'h00;
proc_mem[1159] = 8'h00;
proc_mem[1160] = 8'h00;
proc_mem[1161] = 8'h00;
proc_mem[1162] = 8'h00;
proc_mem[1163] = 8'h00;
proc_mem[1164] = 8'h00;
proc_mem[1165] = 8'h00;
proc_mem[1166] = 8'h00;
proc_mem[1167] = 8'h00;
proc_mem[1168] = 8'h00;
proc_mem[1169] = 8'h00;
proc_mem[1170] = 8'h00;
proc_mem[1171] = 8'h00;
proc_mem[1172] = 8'h00;
proc_mem[1173] = 8'h00;
proc_mem[1174] = 8'h00;
proc_mem[1175] = 8'h00;
proc_mem[1176] = 8'h00;
proc_mem[1177] = 8'h00;
proc_mem[1178] = 8'h00;
proc_mem[1179] = 8'h00;
proc_mem[1180] = 8'h00;
proc_mem[1181] = 8'h00;
proc_mem[1182] = 8'h00;
proc_mem[1183] = 8'h00;
proc_mem[1184] = 8'h00;
proc_mem[1185] = 8'h00;
proc_mem[1186] = 8'h00;
proc_mem[1187] = 8'h00;
proc_mem[1188] = 8'h00;
proc_mem[1189] = 8'h00;
proc_mem[1190] = 8'h00;
proc_mem[1191] = 8'h00;
proc_mem[1192] = 8'h00;
proc_mem[1193] = 8'h00;
proc_mem[1194] = 8'h00;
proc_mem[1195] = 8'h00;
proc_mem[1196] = 8'h00;
proc_mem[1197] = 8'h00;
proc_mem[1198] = 8'h00;
proc_mem[1199] = 8'h00;
proc_mem[1200] = 8'h00;
proc_mem[1201] = 8'h00;
proc_mem[1202] = 8'h00;
proc_mem[1203] = 8'h00;
proc_mem[1204] = 8'h00;
proc_mem[1205] = 8'h00;
proc_mem[1206] = 8'h00;
proc_mem[1207] = 8'h00;
proc_mem[1208] = 8'h00;
proc_mem[1209] = 8'h00;
proc_mem[1210] = 8'h00;
proc_mem[1211] = 8'h00;
proc_mem[1212] = 8'h00;
proc_mem[1213] = 8'h00;
proc_mem[1214] = 8'h00;
proc_mem[1215] = 8'h00;
proc_mem[1216] = 8'h00;
proc_mem[1217] = 8'h00;
proc_mem[1218] = 8'h00;
proc_mem[1219] = 8'h00;
proc_mem[1220] = 8'h00;
proc_mem[1221] = 8'h00;
proc_mem[1222] = 8'h00;
proc_mem[1223] = 8'h00;
proc_mem[1224] = 8'h00;
proc_mem[1225] = 8'h00;
proc_mem[1226] = 8'h00;
proc_mem[1227] = 8'h00;
proc_mem[1228] = 8'h00;
proc_mem[1229] = 8'h00;
proc_mem[1230] = 8'h00;
proc_mem[1231] = 8'h00;
proc_mem[1232] = 8'h00;
proc_mem[1233] = 8'h00;
proc_mem[1234] = 8'h00;
proc_mem[1235] = 8'h00;
proc_mem[1236] = 8'h00;
proc_mem[1237] = 8'h00;
proc_mem[1238] = 8'h00;
proc_mem[1239] = 8'h00;
proc_mem[1240] = 8'h00;
proc_mem[1241] = 8'h00;
proc_mem[1242] = 8'h00;
proc_mem[1243] = 8'h00;
proc_mem[1244] = 8'h00;
proc_mem[1245] = 8'h00;
proc_mem[1246] = 8'h00;
proc_mem[1247] = 8'h00;
proc_mem[1248] = 8'h00;
proc_mem[1249] = 8'h00;
proc_mem[1250] = 8'h00;
proc_mem[1251] = 8'h00;
proc_mem[1252] = 8'h00;
proc_mem[1253] = 8'h00;
proc_mem[1254] = 8'h00;
proc_mem[1255] = 8'h00;
proc_mem[1256] = 8'h00;
proc_mem[1257] = 8'h00;
proc_mem[1258] = 8'h00;
proc_mem[1259] = 8'h00;
proc_mem[1260] = 8'h00;
proc_mem[1261] = 8'h00;
proc_mem[1262] = 8'h00;
proc_mem[1263] = 8'h00;
proc_mem[1264] = 8'h00;
proc_mem[1265] = 8'h00;
proc_mem[1266] = 8'h00;
proc_mem[1267] = 8'h00;
proc_mem[1268] = 8'h00;
proc_mem[1269] = 8'h00;
proc_mem[1270] = 8'h00;
proc_mem[1271] = 8'h00;
proc_mem[1272] = 8'h00;
proc_mem[1273] = 8'h00;
proc_mem[1274] = 8'h00;
proc_mem[1275] = 8'h00;
proc_mem[1276] = 8'h00;
proc_mem[1277] = 8'h00;
proc_mem[1278] = 8'h00;
proc_mem[1279] = 8'h00;
proc_mem[1280] = 8'h00;
proc_mem[1281] = 8'h00;
proc_mem[1282] = 8'h00;
proc_mem[1283] = 8'h00;
proc_mem[1284] = 8'h00;
proc_mem[1285] = 8'h00;
proc_mem[1286] = 8'h00;
proc_mem[1287] = 8'h00;
proc_mem[1288] = 8'h00;
proc_mem[1289] = 8'h00;
proc_mem[1290] = 8'h00;
proc_mem[1291] = 8'h00;
proc_mem[1292] = 8'h00;
proc_mem[1293] = 8'h00;
proc_mem[1294] = 8'h00;
proc_mem[1295] = 8'h00;
proc_mem[1296] = 8'h00;
proc_mem[1297] = 8'h00;
proc_mem[1298] = 8'h00;
proc_mem[1299] = 8'h00;
proc_mem[1300] = 8'h00;
proc_mem[1301] = 8'h00;
proc_mem[1302] = 8'h00;
proc_mem[1303] = 8'h00;
proc_mem[1304] = 8'h00;
proc_mem[1305] = 8'h00;
proc_mem[1306] = 8'h00;
proc_mem[1307] = 8'h00;
proc_mem[1308] = 8'h00;
proc_mem[1309] = 8'h00;
proc_mem[1310] = 8'h00;
proc_mem[1311] = 8'h00;
proc_mem[1312] = 8'h00;
proc_mem[1313] = 8'h00;
proc_mem[1314] = 8'h00;
proc_mem[1315] = 8'h00;
proc_mem[1316] = 8'h00;
proc_mem[1317] = 8'h00;
proc_mem[1318] = 8'h00;
proc_mem[1319] = 8'h00;
proc_mem[1320] = 8'h00;
proc_mem[1321] = 8'h00;
proc_mem[1322] = 8'h00;
proc_mem[1323] = 8'h00;
proc_mem[1324] = 8'h00;
proc_mem[1325] = 8'h00;
proc_mem[1326] = 8'h00;
proc_mem[1327] = 8'h00;
proc_mem[1328] = 8'h00;
proc_mem[1329] = 8'h00;
proc_mem[1330] = 8'h00;
proc_mem[1331] = 8'h00;
proc_mem[1332] = 8'h00;
proc_mem[1333] = 8'h00;
proc_mem[1334] = 8'h00;
proc_mem[1335] = 8'h00;
proc_mem[1336] = 8'h00;
proc_mem[1337] = 8'h00;
proc_mem[1338] = 8'h00;
proc_mem[1339] = 8'h00;
proc_mem[1340] = 8'h00;
proc_mem[1341] = 8'h00;
proc_mem[1342] = 8'h00;
proc_mem[1343] = 8'h00;
proc_mem[1344] = 8'h00;
proc_mem[1345] = 8'h00;
proc_mem[1346] = 8'h00;
proc_mem[1347] = 8'h00;
proc_mem[1348] = 8'h00;
proc_mem[1349] = 8'h00;
proc_mem[1350] = 8'h00;
proc_mem[1351] = 8'h00;
proc_mem[1352] = 8'h00;
proc_mem[1353] = 8'h00;
proc_mem[1354] = 8'h00;
proc_mem[1355] = 8'h00;
proc_mem[1356] = 8'h00;
proc_mem[1357] = 8'h00;
proc_mem[1358] = 8'h00;
proc_mem[1359] = 8'h00;
proc_mem[1360] = 8'h00;
proc_mem[1361] = 8'h00;
proc_mem[1362] = 8'h00;
proc_mem[1363] = 8'h00;
proc_mem[1364] = 8'h00;
proc_mem[1365] = 8'h00;
proc_mem[1366] = 8'h00;
proc_mem[1367] = 8'h00;
proc_mem[1368] = 8'h00;
proc_mem[1369] = 8'h00;
proc_mem[1370] = 8'h00;
proc_mem[1371] = 8'h00;
proc_mem[1372] = 8'h00;
proc_mem[1373] = 8'h00;
proc_mem[1374] = 8'h00;
proc_mem[1375] = 8'h00;
proc_mem[1376] = 8'h00;
proc_mem[1377] = 8'h00;
proc_mem[1378] = 8'h00;
proc_mem[1379] = 8'h00;
proc_mem[1380] = 8'h00;
proc_mem[1381] = 8'h00;
proc_mem[1382] = 8'h00;
proc_mem[1383] = 8'h00;
proc_mem[1384] = 8'h00;
proc_mem[1385] = 8'h00;
proc_mem[1386] = 8'h00;
proc_mem[1387] = 8'h00;
proc_mem[1388] = 8'h00;
proc_mem[1389] = 8'h00;
proc_mem[1390] = 8'h00;
proc_mem[1391] = 8'h00;
proc_mem[1392] = 8'h00;
proc_mem[1393] = 8'h00;
proc_mem[1394] = 8'h00;
proc_mem[1395] = 8'h00;
proc_mem[1396] = 8'h00;
proc_mem[1397] = 8'h00;
proc_mem[1398] = 8'h00;
proc_mem[1399] = 8'h00;
proc_mem[1400] = 8'h00;
proc_mem[1401] = 8'h00;
proc_mem[1402] = 8'h00;
proc_mem[1403] = 8'h00;
proc_mem[1404] = 8'h00;
proc_mem[1405] = 8'h00;
proc_mem[1406] = 8'h00;
proc_mem[1407] = 8'h00;
proc_mem[1408] = 8'h00;
proc_mem[1409] = 8'h00;
proc_mem[1410] = 8'h00;
proc_mem[1411] = 8'h00;
proc_mem[1412] = 8'h00;
proc_mem[1413] = 8'h00;
proc_mem[1414] = 8'h00;
proc_mem[1415] = 8'h00;
proc_mem[1416] = 8'h00;
proc_mem[1417] = 8'h00;
proc_mem[1418] = 8'h00;
proc_mem[1419] = 8'h00;
proc_mem[1420] = 8'h00;
proc_mem[1421] = 8'h00;
proc_mem[1422] = 8'h00;
proc_mem[1423] = 8'h00;
proc_mem[1424] = 8'h00;
proc_mem[1425] = 8'h00;
proc_mem[1426] = 8'h00;
proc_mem[1427] = 8'h00;
proc_mem[1428] = 8'h00;
proc_mem[1429] = 8'h00;
proc_mem[1430] = 8'h00;
proc_mem[1431] = 8'h00;
proc_mem[1432] = 8'h00;
proc_mem[1433] = 8'h00;
proc_mem[1434] = 8'h00;
proc_mem[1435] = 8'h00;
proc_mem[1436] = 8'h00;
proc_mem[1437] = 8'h00;
proc_mem[1438] = 8'h00;
proc_mem[1439] = 8'h00;
proc_mem[1440] = 8'h00;
proc_mem[1441] = 8'h00;
proc_mem[1442] = 8'h00;
proc_mem[1443] = 8'h00;
proc_mem[1444] = 8'h00;
proc_mem[1445] = 8'h00;
proc_mem[1446] = 8'h00;
proc_mem[1447] = 8'h00;
proc_mem[1448] = 8'h00;
proc_mem[1449] = 8'h00;
proc_mem[1450] = 8'h00;
proc_mem[1451] = 8'h00;
proc_mem[1452] = 8'h00;
proc_mem[1453] = 8'h00;
proc_mem[1454] = 8'h00;
proc_mem[1455] = 8'h00;
proc_mem[1456] = 8'h00;
proc_mem[1457] = 8'h00;
proc_mem[1458] = 8'h00;
proc_mem[1459] = 8'h00;
proc_mem[1460] = 8'h00;
proc_mem[1461] = 8'h00;
proc_mem[1462] = 8'h00;
proc_mem[1463] = 8'h00;
proc_mem[1464] = 8'h00;
proc_mem[1465] = 8'h00;
proc_mem[1466] = 8'h00;
proc_mem[1467] = 8'h00;
proc_mem[1468] = 8'h00;
proc_mem[1469] = 8'h00;
proc_mem[1470] = 8'h00;
proc_mem[1471] = 8'h00;
proc_mem[1472] = 8'h00;
proc_mem[1473] = 8'h00;
proc_mem[1474] = 8'h00;
proc_mem[1475] = 8'h00;
proc_mem[1476] = 8'h00;
proc_mem[1477] = 8'h00;
proc_mem[1478] = 8'h00;
proc_mem[1479] = 8'h00;
proc_mem[1480] = 8'h00;
proc_mem[1481] = 8'h00;
proc_mem[1482] = 8'h00;
proc_mem[1483] = 8'h00;
proc_mem[1484] = 8'h00;
proc_mem[1485] = 8'h00;
proc_mem[1486] = 8'h00;
proc_mem[1487] = 8'h00;
proc_mem[1488] = 8'h00;
proc_mem[1489] = 8'h00;
proc_mem[1490] = 8'h00;
proc_mem[1491] = 8'h00;
proc_mem[1492] = 8'h00;
proc_mem[1493] = 8'h00;
proc_mem[1494] = 8'h00;
proc_mem[1495] = 8'h00;
proc_mem[1496] = 8'h00;
proc_mem[1497] = 8'h00;
proc_mem[1498] = 8'h00;
proc_mem[1499] = 8'h00;
proc_mem[1500] = 8'h00;
proc_mem[1501] = 8'h00;
proc_mem[1502] = 8'h00;
proc_mem[1503] = 8'h00;
proc_mem[1504] = 8'h00;
proc_mem[1505] = 8'h00;
proc_mem[1506] = 8'h00;
proc_mem[1507] = 8'h00;
proc_mem[1508] = 8'h00;
proc_mem[1509] = 8'h00;
proc_mem[1510] = 8'h00;
proc_mem[1511] = 8'h00;
proc_mem[1512] = 8'h00;
proc_mem[1513] = 8'h00;
proc_mem[1514] = 8'h00;
proc_mem[1515] = 8'h00;
proc_mem[1516] = 8'h00;
proc_mem[1517] = 8'h00;
proc_mem[1518] = 8'h00;
proc_mem[1519] = 8'h00;
proc_mem[1520] = 8'h00;
proc_mem[1521] = 8'h00;
proc_mem[1522] = 8'h00;
proc_mem[1523] = 8'h00;
proc_mem[1524] = 8'h00;
proc_mem[1525] = 8'h00;
proc_mem[1526] = 8'h00;
proc_mem[1527] = 8'h00;
proc_mem[1528] = 8'h00;
proc_mem[1529] = 8'h00;
proc_mem[1530] = 8'h00;
proc_mem[1531] = 8'h00;
proc_mem[1532] = 8'h00;
proc_mem[1533] = 8'h00;
proc_mem[1534] = 8'h00;
proc_mem[1535] = 8'h00;
proc_mem[1536] = 8'h00;
proc_mem[1537] = 8'h00;
proc_mem[1538] = 8'h00;
proc_mem[1539] = 8'h00;
proc_mem[1540] = 8'h00;
proc_mem[1541] = 8'h00;
proc_mem[1542] = 8'h00;
proc_mem[1543] = 8'h00;
proc_mem[1544] = 8'h00;
proc_mem[1545] = 8'h00;
proc_mem[1546] = 8'h00;
proc_mem[1547] = 8'h00;
proc_mem[1548] = 8'h00;
proc_mem[1549] = 8'h00;
proc_mem[1550] = 8'h00;
proc_mem[1551] = 8'h00;
proc_mem[1552] = 8'h00;
proc_mem[1553] = 8'h00;
proc_mem[1554] = 8'h00;
proc_mem[1555] = 8'h00;
proc_mem[1556] = 8'h00;
proc_mem[1557] = 8'h00;
proc_mem[1558] = 8'h00;
proc_mem[1559] = 8'h00;
proc_mem[1560] = 8'h00;
proc_mem[1561] = 8'h00;
proc_mem[1562] = 8'h00;
proc_mem[1563] = 8'h00;
proc_mem[1564] = 8'h00;
proc_mem[1565] = 8'h00;
proc_mem[1566] = 8'h00;
proc_mem[1567] = 8'h00;
proc_mem[1568] = 8'h00;
proc_mem[1569] = 8'h00;
proc_mem[1570] = 8'h00;
proc_mem[1571] = 8'h00;
proc_mem[1572] = 8'h00;
proc_mem[1573] = 8'h00;
proc_mem[1574] = 8'h00;
proc_mem[1575] = 8'h00;
proc_mem[1576] = 8'h00;
proc_mem[1577] = 8'h00;
proc_mem[1578] = 8'h00;
proc_mem[1579] = 8'h00;
proc_mem[1580] = 8'h00;
proc_mem[1581] = 8'h00;
proc_mem[1582] = 8'h00;
proc_mem[1583] = 8'h00;
proc_mem[1584] = 8'h00;
proc_mem[1585] = 8'h00;
proc_mem[1586] = 8'h00;
proc_mem[1587] = 8'h00;
proc_mem[1588] = 8'h00;
proc_mem[1589] = 8'h00;
proc_mem[1590] = 8'h00;
proc_mem[1591] = 8'h00;
proc_mem[1592] = 8'h00;
proc_mem[1593] = 8'h00;
proc_mem[1594] = 8'h00;
proc_mem[1595] = 8'h00;
proc_mem[1596] = 8'h00;
proc_mem[1597] = 8'h00;
proc_mem[1598] = 8'h00;
proc_mem[1599] = 8'h00;
proc_mem[1600] = 8'h00;
proc_mem[1601] = 8'h00;
proc_mem[1602] = 8'h00;
proc_mem[1603] = 8'h00;
proc_mem[1604] = 8'h00;
proc_mem[1605] = 8'h00;
proc_mem[1606] = 8'h00;
proc_mem[1607] = 8'h00;
proc_mem[1608] = 8'h00;
proc_mem[1609] = 8'h00;
proc_mem[1610] = 8'h00;
proc_mem[1611] = 8'h00;
proc_mem[1612] = 8'h00;
proc_mem[1613] = 8'h00;
proc_mem[1614] = 8'h00;
proc_mem[1615] = 8'h00;
proc_mem[1616] = 8'h00;
proc_mem[1617] = 8'h00;
proc_mem[1618] = 8'h00;
proc_mem[1619] = 8'h00;
proc_mem[1620] = 8'h00;
proc_mem[1621] = 8'h00;
proc_mem[1622] = 8'h00;
proc_mem[1623] = 8'h00;
proc_mem[1624] = 8'h00;
proc_mem[1625] = 8'h00;
proc_mem[1626] = 8'h00;
proc_mem[1627] = 8'h00;
proc_mem[1628] = 8'h00;
proc_mem[1629] = 8'h00;
proc_mem[1630] = 8'h00;
proc_mem[1631] = 8'h00;
proc_mem[1632] = 8'h00;
proc_mem[1633] = 8'h00;
proc_mem[1634] = 8'h00;
proc_mem[1635] = 8'h00;
proc_mem[1636] = 8'h00;
proc_mem[1637] = 8'h00;
proc_mem[1638] = 8'h00;
proc_mem[1639] = 8'h00;
proc_mem[1640] = 8'h00;
proc_mem[1641] = 8'h00;
proc_mem[1642] = 8'h00;
proc_mem[1643] = 8'h00;
proc_mem[1644] = 8'h00;
proc_mem[1645] = 8'h00;
proc_mem[1646] = 8'h00;
proc_mem[1647] = 8'h00;
proc_mem[1648] = 8'h00;
proc_mem[1649] = 8'h00;
proc_mem[1650] = 8'h00;
proc_mem[1651] = 8'h00;
proc_mem[1652] = 8'h00;
proc_mem[1653] = 8'h00;
proc_mem[1654] = 8'h00;
proc_mem[1655] = 8'h00;
proc_mem[1656] = 8'h00;
proc_mem[1657] = 8'h00;
proc_mem[1658] = 8'h00;
proc_mem[1659] = 8'h00;
proc_mem[1660] = 8'h00;
proc_mem[1661] = 8'h00;
proc_mem[1662] = 8'h00;
proc_mem[1663] = 8'h00;
proc_mem[1664] = 8'h00;
proc_mem[1665] = 8'h00;
proc_mem[1666] = 8'h00;
proc_mem[1667] = 8'h00;
proc_mem[1668] = 8'h00;
proc_mem[1669] = 8'h00;
proc_mem[1670] = 8'h00;
proc_mem[1671] = 8'h00;
proc_mem[1672] = 8'h00;
proc_mem[1673] = 8'h00;
proc_mem[1674] = 8'h00;
proc_mem[1675] = 8'h00;
proc_mem[1676] = 8'h00;
proc_mem[1677] = 8'h00;
proc_mem[1678] = 8'h00;
proc_mem[1679] = 8'h00;
proc_mem[1680] = 8'h00;
proc_mem[1681] = 8'h00;
proc_mem[1682] = 8'h00;
proc_mem[1683] = 8'h00;
proc_mem[1684] = 8'h00;
proc_mem[1685] = 8'h00;
proc_mem[1686] = 8'h00;
proc_mem[1687] = 8'h00;
proc_mem[1688] = 8'h00;
proc_mem[1689] = 8'h00;
proc_mem[1690] = 8'h00;
proc_mem[1691] = 8'h00;
proc_mem[1692] = 8'h00;
proc_mem[1693] = 8'h00;
proc_mem[1694] = 8'h00;
proc_mem[1695] = 8'h00;
proc_mem[1696] = 8'h00;
proc_mem[1697] = 8'h00;
proc_mem[1698] = 8'h00;
proc_mem[1699] = 8'h00;
proc_mem[1700] = 8'h00;
proc_mem[1701] = 8'h00;
proc_mem[1702] = 8'h00;
proc_mem[1703] = 8'h00;
proc_mem[1704] = 8'h00;
proc_mem[1705] = 8'h00;
proc_mem[1706] = 8'h00;
proc_mem[1707] = 8'h00;
proc_mem[1708] = 8'h00;
proc_mem[1709] = 8'h00;
proc_mem[1710] = 8'h00;
proc_mem[1711] = 8'h00;
proc_mem[1712] = 8'h00;
proc_mem[1713] = 8'h00;
proc_mem[1714] = 8'h00;
proc_mem[1715] = 8'h00;
proc_mem[1716] = 8'h00;
proc_mem[1717] = 8'h00;
proc_mem[1718] = 8'h00;
proc_mem[1719] = 8'h00;
proc_mem[1720] = 8'h00;
proc_mem[1721] = 8'h00;
proc_mem[1722] = 8'h00;
proc_mem[1723] = 8'h00;
proc_mem[1724] = 8'h00;
proc_mem[1725] = 8'h00;
proc_mem[1726] = 8'h00;
proc_mem[1727] = 8'h00;
proc_mem[1728] = 8'h00;
proc_mem[1729] = 8'h00;
proc_mem[1730] = 8'h00;
proc_mem[1731] = 8'h00;
proc_mem[1732] = 8'h00;
proc_mem[1733] = 8'h00;
proc_mem[1734] = 8'h00;
proc_mem[1735] = 8'h00;
proc_mem[1736] = 8'h00;
proc_mem[1737] = 8'h00;
proc_mem[1738] = 8'h00;
proc_mem[1739] = 8'h00;
proc_mem[1740] = 8'h00;
proc_mem[1741] = 8'h00;
proc_mem[1742] = 8'h00;
proc_mem[1743] = 8'h00;
proc_mem[1744] = 8'h00;
proc_mem[1745] = 8'h00;
proc_mem[1746] = 8'h00;
proc_mem[1747] = 8'h00;
proc_mem[1748] = 8'h00;
proc_mem[1749] = 8'h00;
proc_mem[1750] = 8'h00;
proc_mem[1751] = 8'h00;
proc_mem[1752] = 8'h00;
proc_mem[1753] = 8'h00;
proc_mem[1754] = 8'h00;
proc_mem[1755] = 8'h00;
proc_mem[1756] = 8'h00;
proc_mem[1757] = 8'h00;
proc_mem[1758] = 8'h00;
proc_mem[1759] = 8'h00;
proc_mem[1760] = 8'h00;
proc_mem[1761] = 8'h00;
proc_mem[1762] = 8'h00;
proc_mem[1763] = 8'h00;
proc_mem[1764] = 8'h00;
proc_mem[1765] = 8'h00;
proc_mem[1766] = 8'h00;
proc_mem[1767] = 8'h00;
proc_mem[1768] = 8'h00;
proc_mem[1769] = 8'h00;
proc_mem[1770] = 8'h00;
proc_mem[1771] = 8'h00;
proc_mem[1772] = 8'h00;
proc_mem[1773] = 8'h00;
proc_mem[1774] = 8'h00;
proc_mem[1775] = 8'h00;
proc_mem[1776] = 8'h00;
proc_mem[1777] = 8'h00;
proc_mem[1778] = 8'h00;
proc_mem[1779] = 8'h00;
proc_mem[1780] = 8'h00;
proc_mem[1781] = 8'h00;
proc_mem[1782] = 8'h00;
proc_mem[1783] = 8'h00;
proc_mem[1784] = 8'h00;
proc_mem[1785] = 8'h00;
proc_mem[1786] = 8'h00;
proc_mem[1787] = 8'h00;
proc_mem[1788] = 8'h00;
proc_mem[1789] = 8'h00;
proc_mem[1790] = 8'h00;
proc_mem[1791] = 8'h00;
proc_mem[1792] = 8'h00;
proc_mem[1793] = 8'h00;
proc_mem[1794] = 8'h00;
proc_mem[1795] = 8'h00;
proc_mem[1796] = 8'h00;
proc_mem[1797] = 8'h00;
proc_mem[1798] = 8'h00;
proc_mem[1799] = 8'h00;
proc_mem[1800] = 8'h00;
proc_mem[1801] = 8'h00;
proc_mem[1802] = 8'h00;
proc_mem[1803] = 8'h00;
proc_mem[1804] = 8'h00;
proc_mem[1805] = 8'h00;
proc_mem[1806] = 8'h00;
proc_mem[1807] = 8'h00;
proc_mem[1808] = 8'h00;
proc_mem[1809] = 8'h00;
proc_mem[1810] = 8'h00;
proc_mem[1811] = 8'h00;
proc_mem[1812] = 8'h00;
proc_mem[1813] = 8'h00;
proc_mem[1814] = 8'h00;
proc_mem[1815] = 8'h00;
proc_mem[1816] = 8'h00;
proc_mem[1817] = 8'h00;
proc_mem[1818] = 8'h00;
proc_mem[1819] = 8'h00;
proc_mem[1820] = 8'h00;
proc_mem[1821] = 8'h00;
proc_mem[1822] = 8'h00;
proc_mem[1823] = 8'h00;
proc_mem[1824] = 8'h00;
proc_mem[1825] = 8'h00;
proc_mem[1826] = 8'h00;
proc_mem[1827] = 8'h00;
proc_mem[1828] = 8'h00;
proc_mem[1829] = 8'h00;
proc_mem[1830] = 8'h00;
proc_mem[1831] = 8'h00;
proc_mem[1832] = 8'h00;
proc_mem[1833] = 8'h00;
proc_mem[1834] = 8'h00;
proc_mem[1835] = 8'h00;
proc_mem[1836] = 8'h00;
proc_mem[1837] = 8'h00;
proc_mem[1838] = 8'h00;
proc_mem[1839] = 8'h00;
proc_mem[1840] = 8'h00;
proc_mem[1841] = 8'h00;
proc_mem[1842] = 8'h00;
proc_mem[1843] = 8'h00;
proc_mem[1844] = 8'h00;
proc_mem[1845] = 8'h00;
proc_mem[1846] = 8'h00;
proc_mem[1847] = 8'h00;
proc_mem[1848] = 8'h00;
proc_mem[1849] = 8'h00;
proc_mem[1850] = 8'h00;
proc_mem[1851] = 8'h00;
proc_mem[1852] = 8'h00;
proc_mem[1853] = 8'h00;
proc_mem[1854] = 8'h00;
proc_mem[1855] = 8'h00;
proc_mem[1856] = 8'h00;
proc_mem[1857] = 8'h00;
proc_mem[1858] = 8'h00;
proc_mem[1859] = 8'h00;
proc_mem[1860] = 8'h00;
proc_mem[1861] = 8'h00;
proc_mem[1862] = 8'h00;
proc_mem[1863] = 8'h00;
proc_mem[1864] = 8'h00;
proc_mem[1865] = 8'h00;
proc_mem[1866] = 8'h00;
proc_mem[1867] = 8'h00;
proc_mem[1868] = 8'h00;
proc_mem[1869] = 8'h00;
proc_mem[1870] = 8'h00;
proc_mem[1871] = 8'h00;
proc_mem[1872] = 8'h00;
proc_mem[1873] = 8'h00;
proc_mem[1874] = 8'h00;
proc_mem[1875] = 8'h00;
proc_mem[1876] = 8'h00;
proc_mem[1877] = 8'h00;
proc_mem[1878] = 8'h00;
proc_mem[1879] = 8'h00;
proc_mem[1880] = 8'h00;
proc_mem[1881] = 8'h00;
proc_mem[1882] = 8'h00;
proc_mem[1883] = 8'h00;
proc_mem[1884] = 8'h00;
proc_mem[1885] = 8'h00;
proc_mem[1886] = 8'h00;
proc_mem[1887] = 8'h00;
proc_mem[1888] = 8'h00;
proc_mem[1889] = 8'h00;
proc_mem[1890] = 8'h00;
proc_mem[1891] = 8'h00;
proc_mem[1892] = 8'h00;
proc_mem[1893] = 8'h00;
proc_mem[1894] = 8'h00;
proc_mem[1895] = 8'h00;
proc_mem[1896] = 8'h00;
proc_mem[1897] = 8'h00;
proc_mem[1898] = 8'h00;
proc_mem[1899] = 8'h00;
proc_mem[1900] = 8'h00;
proc_mem[1901] = 8'h00;
proc_mem[1902] = 8'h00;
proc_mem[1903] = 8'h00;
proc_mem[1904] = 8'h00;
proc_mem[1905] = 8'h00;
proc_mem[1906] = 8'h00;
proc_mem[1907] = 8'h00;
proc_mem[1908] = 8'h00;
proc_mem[1909] = 8'h00;
proc_mem[1910] = 8'h00;
proc_mem[1911] = 8'h00;
proc_mem[1912] = 8'h00;
proc_mem[1913] = 8'h00;
proc_mem[1914] = 8'h00;
proc_mem[1915] = 8'h00;
proc_mem[1916] = 8'h00;
proc_mem[1917] = 8'h00;
proc_mem[1918] = 8'h00;
proc_mem[1919] = 8'h00;
proc_mem[1920] = 8'h00;
proc_mem[1921] = 8'h00;
proc_mem[1922] = 8'h00;
proc_mem[1923] = 8'h00;
proc_mem[1924] = 8'h00;
proc_mem[1925] = 8'h00;
proc_mem[1926] = 8'h00;
proc_mem[1927] = 8'h00;
proc_mem[1928] = 8'h00;
proc_mem[1929] = 8'h00;
proc_mem[1930] = 8'h00;
proc_mem[1931] = 8'h00;
proc_mem[1932] = 8'h00;
proc_mem[1933] = 8'h00;
proc_mem[1934] = 8'h00;
proc_mem[1935] = 8'h00;
proc_mem[1936] = 8'h00;
proc_mem[1937] = 8'h00;
proc_mem[1938] = 8'h00;
proc_mem[1939] = 8'h00;
proc_mem[1940] = 8'h00;
proc_mem[1941] = 8'h00;
proc_mem[1942] = 8'h00;
proc_mem[1943] = 8'h00;
proc_mem[1944] = 8'h00;
proc_mem[1945] = 8'h00;
proc_mem[1946] = 8'h00;
proc_mem[1947] = 8'h00;
proc_mem[1948] = 8'h00;
proc_mem[1949] = 8'h00;
proc_mem[1950] = 8'h00;
proc_mem[1951] = 8'h00;
proc_mem[1952] = 8'h00;
proc_mem[1953] = 8'h00;
proc_mem[1954] = 8'h00;
proc_mem[1955] = 8'h00;
proc_mem[1956] = 8'h00;
proc_mem[1957] = 8'h00;
proc_mem[1958] = 8'h00;
proc_mem[1959] = 8'h00;
proc_mem[1960] = 8'h00;
proc_mem[1961] = 8'h00;
proc_mem[1962] = 8'h00;
proc_mem[1963] = 8'h00;
proc_mem[1964] = 8'h00;
proc_mem[1965] = 8'h00;
proc_mem[1966] = 8'h00;
proc_mem[1967] = 8'h00;
proc_mem[1968] = 8'h00;
proc_mem[1969] = 8'h00;
proc_mem[1970] = 8'h00;
proc_mem[1971] = 8'h00;
proc_mem[1972] = 8'h00;
proc_mem[1973] = 8'h00;
proc_mem[1974] = 8'h00;
proc_mem[1975] = 8'h00;
proc_mem[1976] = 8'h00;
proc_mem[1977] = 8'h00;
proc_mem[1978] = 8'h00;
proc_mem[1979] = 8'h00;
proc_mem[1980] = 8'h00;
proc_mem[1981] = 8'h00;
proc_mem[1982] = 8'h00;
proc_mem[1983] = 8'h00;
proc_mem[1984] = 8'h00;
proc_mem[1985] = 8'h00;
proc_mem[1986] = 8'h00;
proc_mem[1987] = 8'h00;
proc_mem[1988] = 8'h00;
proc_mem[1989] = 8'h00;
proc_mem[1990] = 8'h00;
proc_mem[1991] = 8'h00;
proc_mem[1992] = 8'h00;
proc_mem[1993] = 8'h00;
proc_mem[1994] = 8'h00;
proc_mem[1995] = 8'h00;
proc_mem[1996] = 8'h00;
proc_mem[1997] = 8'h00;
proc_mem[1998] = 8'h00;
proc_mem[1999] = 8'h00;
proc_mem[2000] = 8'h00;
proc_mem[2001] = 8'h00;
proc_mem[2002] = 8'h00;
proc_mem[2003] = 8'h00;
proc_mem[2004] = 8'h00;
proc_mem[2005] = 8'h00;
proc_mem[2006] = 8'h00;
proc_mem[2007] = 8'h00;
proc_mem[2008] = 8'h00;
proc_mem[2009] = 8'h00;
proc_mem[2010] = 8'h00;
proc_mem[2011] = 8'h00;
proc_mem[2012] = 8'h00;
proc_mem[2013] = 8'h00;
proc_mem[2014] = 8'h00;
proc_mem[2015] = 8'h00;
proc_mem[2016] = 8'h00;
proc_mem[2017] = 8'h00;
proc_mem[2018] = 8'h00;
proc_mem[2019] = 8'h00;
proc_mem[2020] = 8'h00;
proc_mem[2021] = 8'h00;
proc_mem[2022] = 8'h00;
proc_mem[2023] = 8'h00;
proc_mem[2024] = 8'h00;
proc_mem[2025] = 8'h00;
proc_mem[2026] = 8'h00;
proc_mem[2027] = 8'h00;
proc_mem[2028] = 8'h00;
proc_mem[2029] = 8'h00;
proc_mem[2030] = 8'h00;
proc_mem[2031] = 8'h00;
proc_mem[2032] = 8'h00;
proc_mem[2033] = 8'h00;
proc_mem[2034] = 8'h00;
proc_mem[2035] = 8'h00;
proc_mem[2036] = 8'h00;
proc_mem[2037] = 8'h00;
proc_mem[2038] = 8'h00;
proc_mem[2039] = 8'h00;
proc_mem[2040] = 8'h00;
proc_mem[2041] = 8'h00;
proc_mem[2042] = 8'h00;
proc_mem[2043] = 8'h00;
proc_mem[2044] = 8'h00;
proc_mem[2045] = 8'h00;
proc_mem[2046] = 8'h00;
proc_mem[2047] = 8'h00;

		
		
		//proc_mem[4095] = 8'b0;
		//proc_mem[0] = 8'h
		//proc_mem[0] = 8'h
		//proc_mem[0] = 8'h
		//proc_mem[0] = 8'h
		//proc_mem[0] = 8'h
		//proc_mem[0] = 8'h
		//proc_mem[0] = 8'h
		//proc_mem[0] = 8'h
		//proc_mem[0] = 8'h
		//proc_mem[0] = 8'h
		//proc_mem[0] = 8'h
		//proc_mem[0] = 8'h
		//proc_mem[0] = 8'h
		//proc_mem[0] = 8'h
		
		
	end
	
	always@(*)
	begin
		
		imem_error=0;
		if(PC>4095)
		begin
			imem_error=1;
		end
		
		
		
		instr = {
			proc_mem[PC],
			proc_mem[PC+1],
			proc_mem[PC+2],
			proc_mem[PC+3],
			proc_mem[PC+4],
			proc_mem[PC+5],
			proc_mem[PC+6],
			proc_mem[PC+7],
			proc_mem[PC+8],
			proc_mem[PC+9]
			};
		
		instr2 = {
			proc_mem[PC+9],
			proc_mem[PC+8],
			proc_mem[PC+7],
			proc_mem[PC+6],
			proc_mem[PC+5],
			proc_mem[PC+4],
			proc_mem[PC+3],
			proc_mem[PC+2],
			proc_mem[PC+1],
			proc_mem[PC]
			};
				
			
		$display("instr=%x", instr);
		
		icode = instr[0:3]; // high nibble
		ifun = instr[4:7]; //low nibble
		
		instr_validity = 1'b1;
		
		// go through all icode cases
		// halt 0x00
		if(icode==4'b0000)
		begin
			hlt=1;
			valP = PC+64'd1;
		end
		// nop 0x10
		else if(icode==4'b0001)
		begin
			valP = PC+64'd1;
		end
		// cmovxx 0x2Fn
		else if(icode==4'b0010)
		begin
			rA = instr[8:11]; // register number
			rB = instr[12:15]; // register number
			valP = PC+64'd2;
		end
		// irmov 0x30
		else if(icode==4'b0011)
		begin
			rA = instr[8:11]; // register number
			rB = instr[12:15]; // register number
			valC = instr2[79:16];
			valP = PC+64'd10;
		end
		// rmmov 0x40
		else if(icode==4'b0100)
		begin
			rA = instr[8:11]; // register number
			rB = instr[12:15]; // register number
			valC = instr2[79:16];
			valP = PC+64'd10;
		end
		// mrmov 0x50
		else if(icode==4'b0101)
		begin
			rA = instr[8:11]; // register number
			rB = instr[12:15]; // register number
			valC = instr2[79:16];
			valP = PC+64'd10;
		end
		// OP 0x6Fn	
		else if(icode==4'b0110)
		begin
			rA = instr[8:11]; // register number
			rB = instr[12:15]; // register number
			valP = PC+64'd2;
		end
		// jXX 0x7Fn	
		else if(icode==4'b0111)
		begin
			valC = instr2[71:8];
			valP = PC+64'd9;
		end
		// call 0x80
		else if(icode==4'b1000)
		begin
			valC = instr2[71:8];
			valP = instr[8:15];//PC+64'd9;
		end
		// ret 0x90	
		else if(icode==4'b1001)
		begin
			valP = PC+64'd1;
		end
		// pushq 0xa0	
		else if(icode==4'b1010)
		begin
			rA = instr[8:11]; // register number
			rB = instr[12:15]; // register number
			valP = PC+64'd2;
		end
		// popq 0xb0	
		else if(icode==4'b1011)
		begin
			rA = instr[8:11]; // register number
			rB = instr[12:15]; // register number
			valP = PC+64'd2;
		end
		else begin
			instr_validity=1'b0;
		end
		
		$display("rA=%d, rB=%d, valC=%x, valP=%d", rA, rB, valC, valP);
		
	
	
	end
	
	endmodule
	